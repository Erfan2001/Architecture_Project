`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:41:36 06/24/2021 
// Design Name: 
// Module Name:    ALU_CTR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU_CTR(
		input [5:0]func,
		input [5:0] opcode,
		output [2:0] alu_op
    );
	 
	 


endmodule
