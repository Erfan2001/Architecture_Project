`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:34:29 06/26/2021 
// Design Name: 
// Module Name:    Jump_Mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Jump_Mux(
		input [31:0] zero_base,
		input branch,
		output [31:0] resultMuxFromMem
    );
	always@(*)
		begin
			
		end

endmodule
